module PE(
	input clk,
	input rst,
	input SPIKE_in0,
	input SPIKE_in1,
	input SPIKE_in2,
	input SPIKE_in3,
	input [7:0] WEIGHT_IN,
	input EN,
	input layer,
	output SPIKE_OUT
);


endmodule